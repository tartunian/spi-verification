`define HALF_CLK_PRD	10